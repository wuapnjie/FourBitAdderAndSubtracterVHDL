----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:31:48 05/17/2016 
-- Design Name: 
-- Module Name:    TwoBitAdder - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity OneBitAdder is
    Port ( 
			  A : in  STD_LOGIC;
           B : in  STD_LOGIC;
           Cin : in  STD_LOGIC;
           O : out  STD_LOGIC;
           Cout : out  STD_LOGIC);
end OneBitAdder;

architecture Behavioral of OneBitAdder is

begin
	O<=A xor B xor Cin;
	Cout <= (A and Cin) or (B and Cin) or (A and B);

end Behavioral;